../isat_calc_v1_0/iSat.vhd